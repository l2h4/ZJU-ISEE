.SUBCKT OPAMP 1 11 14 15 2 6
*1  VDD
*11 VSS
*14 Vip
*15 Vin
*2  Vop
*6  Von

M1 8 14 13 13 p08 W=300u L=3u
M2 9 15 13 13 p08 W=300u L=3u
M3 13 12 1 1 p08 W=600u L=3u
M4 3 2 1 1 p08 W=360u L=3u
M5 4 2 1 1 p08 W=360u L=3u
M6 2 5 3 3 p08 W=360u L=3u
M7 6 5 4 4 p08 W=360u L=3u
M8 2 7 8 8 n08 W=280u L=4u
M9 6 7 9 9 n08 W=280u L=4u
M10 8 10 11 11 n08 W=280u L=4u
M11 9 10 11 11 n08 W=280u L=4u
M12 16 12 1 1 p08 W=28u L=4u
M13 18 10 11 11 n08 W=12u L=4u
M14 10 7 18 18 n08 W=12u L=4u
M15 12 5 16 16 p08 W=28u L=4u
M16 17 12 1 1 p08 W=28u L=4u
M17 7 5 17 17 p08 W=28u L=4u
R0 12 5 35K
R1 7 10 50K
IBIAS 5 11 10u


.MODEL n08 NMOS VTO = 0.70 KP = 110U GAMMA = 0.4  LAMBDA = 0.04 
+ PHI = 0.7 MJ = 0.5 MJSW = 0.38 CGBO = 700P CGSO = 220P CGDO = 220P 
+ CJ = 770U CJSW = 380P LD = 0.016U TOX = 14N
.MODEL p08 PMOS VTO = -0.70 KP = 50U GAMMA = 0.57 LAMBDA = 0.05 
+ PHI = 0.8 MJ = 0.5 MJSW = 0.35 CGBO = 700P CGSO = 220P CGDO = 220P 
+ CJ = 560U CJSW = 350P LD = 0.014U TOX = 14N

.ENDS