.SUBCKT SWITCH 2 3 7 10 12
* 2 vin
* 3 vout
* 7 vclk
* 10 VDD
* 12 vclkf
M1 3 1 2 0 n08 W=714u L=1u 
M2 1 4 5 5 p08 W=89u L=1u
M3 2 1 6 0 n08 W=178u L=1u
M4 9 7 0 0 n08 W=357u L=1u
M5 5 1 10 5 p08 W=178u L=1u
M6 6 7 0 0 n08 W=89u L=1u
M8 1 10 9 0 n08 W=357u L=1u
Ma 4 12 6 0 n08 W=9u L=1u
Mb 4 12 10 0 p08 W=36 L=1u
Mc 4 1 6 0 n08 W=178u L=1u
C1 3 8 0.5p
CB 5 6 0.25p

.MODEL n08 NMOS VTO = 0.70 KP = 110U GAMMA = 0.4  LAMBDA = 0.04 
+ PHI = 0.7 MJ = 0.5 MJSW = 0.38 CGBO = 700P CGSO = 220P CGDO = 220P 
+ CJ = 770U CJSW = 380P LD = 0.016U TOX = 14N
.MODEL p08 PMOS VTO = -0.70 KP = 50U GAMMA = 0.57 LAMBDA = 0.05 
+ PHI = 0.8 MJ = 0.5 MJSW = 0.35 CGBO = 700P CGSO = 220P CGDO = 220P 
+ CJ = 560U CJSW = 350P LD = 0.014U TOX = 14N

.ENDS