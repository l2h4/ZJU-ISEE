.SUBCKT OPAMP 1 2 7 8 10 11
*1 vin
*2 vip
*7 VDD
*8 VSS
*10 vop
*11 von
M1 3 1 5 5 n08 W=8u L=1u
M2 4 2 5 5 n08 W=8u L=1u
M3 3 4 7 7 p08 W=23u L=1u
M4 4 4 7 7 p08 W=23u L=1u
M5 5 9 8 8 n08 W=4u L=1u
M6 11 4 7 7 p08 W=190u L=1u
M7 11 9 8 8 n08 W=17u L=1u
M8 9 9 8 8 n08 W=4u L=1u
M9 10 9 8 8 n08 W=17u L=1u
M10 10 3 7 7 p08 W=190u L=1u
C1 4 11 3p
C2 3 10 3p
IBIA 7 9 30U

.MODEL n08 NMOS VTO = 0.70 KP = 110U GAMMA = 0.4  LAMBDA = 0.04 
+ PHI = 0.7 MJ = 0.5 MJSW = 0.38 CGBO = 700P CGSO = 220P CGDO = 220P 
+ CJ = 770U CJSW = 380P LD = 0.016U TOX = 14N
.MODEL p08 PMOS VTO = -0.70 KP = 50U GAMMA = 0.57 LAMBDA = 0.05 
+ PHI = 0.8 MJ = 0.5 MJSW = 0.35 CGBO = 700P CGSO = 220P CGDO = 220P 
+ CJ = 560U CJSW = 350P LD = 0.014U TOX = 14N

.ENDS
