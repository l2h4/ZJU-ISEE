.title OPA_CMRR

.include 'OPA.cdl'

x1 1 2 3 4 5 6 OPAMP
*1 vin
*2 vip
*3 VDD
*4 VSS
*5 vop
*6 von
VDD 3 0 DC  5
VSS 0 4 DC  5
C1 5 0 10P
C2 6 0 10p
.PARAM VCM=1
VCM1 1 0 DC 0 AC VCM
VCM2 2 6 DC 0 AC VCM 

.ac dec 10 1 1g
.probe ac vdb(6) vp(6)
.probe ac cmrr_db=par('- vdb(6)') cmrr_phase=par('- vp(6)')

.temp 27								
.option post accurate probe

.end